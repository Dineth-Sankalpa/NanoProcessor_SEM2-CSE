library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity NanoProcessor_Sim is
--  Port ( );
end NanoProcessor_Sim;

architecture Behavioral of NanoProcessor_Sim is

component NanoProcessor_Nano4ce
     Port ( 
        Clk               : in  STD_LOGIC;
        Reset             : in  STD_LOGIC;
        
        Zero_Flag_LED     : out STD_LOGIC;
        Overflow_Flag_LED : out STD_LOGIC;
        Jump_Flag_LED     : out STD_LOGIC;
        NEG_FLAG_LED      : out STD_LOGIC;
        
        R7_Out            : out STD_LOGIC_VECTOR(3 downto 0);
        sevenSeg          : out STD_LOGIC_VECTOR(6 downto 0);
        Display           : out STD_LOGIC_VECTOR(3 downto 0);
        SW14, SW15              : in STD_LOGIC
    );
end component;

signal Clk, Reset, Zero_Flag_LED, Overflow_Flag_LED, Jump_Flag_LED, NEG_FLAG_LED  : std_logic;
signal R7_Out, Display : STD_LOGIC_VECTOR(3 downto 0);
signal sevenSeg : STD_LOGIC_VECTOR(6 downto 0);
signal sw14_tb: std_logic := '0';  -- Or whatever initial value you want
signal sw15_tb: std_logic := '0';  -- Or whatever initial value you want

begin

UUT: NanoProcessor_Nano4ce
    port map (
        Clk                => Clk,
        Reset              => Reset,
        Zero_Flag_LED      => Zero_Flag_LED,
        Overflow_Flag_LED  => Overflow_Flag_LED,
        Jump_Flag_LED      => Jump_Flag_LED,
        NEG_FLAG_LED       => NEG_FLAG_LED,
        R7_Out             => R7_Out,
        sevenSeg           => sevenSeg,
        Display            => Display,
        SW14               => sw14_tb,
        SW15               => sw15_tb
);

clk_process : process
begin
    Clk <= '0';
    wait for 10ns;
    
    Clk <= '1';
    wait for 10ns;
end process;

--Process_Sim : process
--begin



end Behavioral;