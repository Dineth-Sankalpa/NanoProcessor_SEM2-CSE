library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL; -- for arithmetic functions

entity LUT_16_7 is
    Port ( 
        address_LUT : in STD_LOGIC_VECTOR (3 downto 0);
        data_LUT : out STD_LOGIC_VECTOR (6 downto 0)
    );
end LUT_16_7;

architecture Behavioral of LUT_16_7 is
    type rom_type is array (0 to 15) of std_logic_vector(6 downto 0);
    
    signal sevenSegment_ROM : rom_type := (
        "1000000", -- 0
        "1111001", -- 1
        "0100100", -- 2
        "0110000", -- 3
        "0011001", -- 4
        "0010010", -- 5
        "0000010", -- 6
        "1111000", -- 7
        "0000000", -- 8
        "0010000", -- 9
        "0001000", -- a
        "0000011", -- b
        "1000110", -- c
        "0100001", -- d
        "0000110", -- e
--        "0001110"  -- f
        "0111111"  -- '-'
   );

begin
    process(address_LUT)
        begin
            data_LUT <= sevenSegment_ROM(to_integer(unsigned(address_LUT)));
    end process;

end Behavioral;
